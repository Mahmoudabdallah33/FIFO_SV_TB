
//import pkg::*;
interface dut_if ();

bit clk1,clk2; logic rst, wrt, rd;
logic [31:0] data_in;
logic [31:0] data_out;






endinterface
