package pkg_1;
typedef class transaction;
typedef class generator;
typedef class driver;
typedef class monitor_in;
typedef class check;
typedef class env;


`include"transaction.sv"
`include"generator.sv"
`include"driver.sv"
`include"monitor_in.sv"
`include"checker.sv"
`include"enviroment.sv"


endpackage
